--| Nhóm                | Thủ tục / Hàm                                                                                         | Nhiệm vụ                                                                      | Khi dùng                                        |
--| ------------------- | ----------------------------------------------------------------------------------------------------- | ----------------------------------------------------------------------------- | ----------------------------------------------- |
--| **Khởi tạo**        | `NewID`                                                                                               | Tạo **CoverageID**, gieo seed ngẫu nhiên                                      | Trước khi AddBins/ICover                        |
--| **Mô hình (Item)**  | `GenBin`, `IllegalBin`, `IgnoreBin` → `AddBins`                                                       | Khai báo các **bin** giá trị / phạm vi                                        | Theo test‑plan item coverage                    |
--| **Mô hình (Cross)** | `AddCross` + nhiều `GenBin`                                                                           | Tạo ma trận quan hệ (đến 20 item)                                             | Kiểm tra tổ hợp thanh ghi, cổng…                |
--| **Tích lũy**        | `ICover`                                                                                              | Ghi giá trị (int / int\_vector) vào mô hình                                   | Clock‑sampling, transaction‑sampling            |
--| **Kết thúc?**       | `IsCovered`                                                                                           | TRUE khi mọi bin đạt goal                                                     | Dừng test nhanh                                 |
--| **Thống kê**        | `GetCov`, `GetItemCount`, `GetTotalCovGoal`                                                           | % cover, số mục đã lấy                                                        | Báo cáo CI                                      |
--| **Random hóc cao**  | `GetRandPoint`, `GetRandBinVal`                                                                       | “Intelligent Coverage” bốc **lỗ hổng**                                        | Giảm mô phỏng từ N·logN xuống ≈ N turn1file17 |
--| **Báo cáo**         | `WriteBin`, `WriteCovHoles`, `FileOpenWriteBin`                                                       | Xuất bảng bin hoặc chỉ “hole”                                                 | Thân thiện requirements tools                   |
--| **Điều khiển**      | `SetIllegalMode`, `SetBinSize`, `SetWeightMode`, `SetCovTarget`, `SetCovThreshold`, `SetCountMode`, … | Tắt ALERT cho bin illegal, tối ưu RAM, chỉnh trọng số random, đặt ngưỡng %... | Nâng cao / tối ưu turn1file9                  |
--| **Transition**      | `TCover`                                                                                              | Bao phủ **chuỗi** giá trị                                                     | FSM, giao thức handshake                        |
--| **Tiện ích**        | `IsInitialized`, `GetSeed`, `SetSeed`, `GetRandIndex`, …                                              | Kiểm tra mô hình, tái lập bug                                                 | Debug, regression                               |




library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library OSVVM;
context OSVVM.OSVVMContext;
use osvvm.ScoreboardPkg_slv.all;

entity Test23_Coverage is
end entity;

architecture tb of Test23_Coverage is

constant TB_ID : AlertLogIDType := NewID("Test23_Coverage");
constant SB_ID : ScoreboardIdType := NewID("Scoreboard", TB_ID);
constant COV_ID: CoverageIdType := NewID("Coverage", TB_ID);


begin

    Test_proc: process
    begin

        SetTestName("Test23_Coverage");
        SetLogEnable(TB_ID,PASSED, TRUE);
        SetLogEnable(TB_ID,INFO, TRUE);
        TranscriptOpen;
        SetTranscriptMirror(TRUE);

        wait for 0 ns; wait for 0 ns;
        AddBins(COV_ID, GenBin(1, 3)); -- 3 bin 1, 2, 3
        AddBins(COV_ID, GenBin(4,252,2));
        AddBins(COV_ID, GenBin(253, 255));
        wait for 10 ns;

        for i in 0 to 300 loop
            ICover(COV_ID, i);
            Log(TB_ID, "i = " & to_string(i), INFO);
            exit when IsCovered(COV_ID);
        end loop;
        
        wait for 10 ns;
        AffirmIfEqual(TB_ID, IsCovered(COV_ID), TRUE, "Coverage is 100%");
        WriteBin(COV_ID);
        WriteCovHoles(COV_ID); -- in ra hole rong -> neu khong co hole thi khong in ra
        TranscriptClose;
        EndOfTestSummary(ReportAll => TRUE);

        std.env.stop;

    end process;
    
end architecture;